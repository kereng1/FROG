module memory_tb;

  // ============================
  // Parameters
  // ============================
  localparam IMEM_SIZE_WORDS = 256;
  localparam DMEM_SIZE_BYTES = 1024;

  // ============================
  // Clock / Reset
  // ============================
  logic clk;
  logic rst;

  always #5 clk = ~clk;

  // ============================
  // DUT signals
  // ============================
  logic [31:0] pc_Q100H;
  logic        ready_Q101H;
  logic [31:0] instruction_Q101H;

  logic [31:0] alu_out_Q103H;
  logic [31:0] dmem_wr_data_Q103H;
  logic        dmem_wr_en_Q103H;
  logic [3:0]  dmem_byte_en_Q103H;
  logic        dmem_is_signed_Q103H;
  logic [31:0] dmem_rd_data_Q104H;

  // ============================
  // DUT instantiation
  // ============================
  memory #(
    .IMEM_SIZE_WORDS(IMEM_SIZE_WORDS),
    .DMEM_SIZE_BYTES(DMEM_SIZE_BYTES)
  ) dut (
    .clk(clk),
    .rst(rst),

    .pc_Q100H(pc_Q100H),
    .ready_Q101H(ready_Q101H),
    .instruction_Q101H(instruction_Q101H),

    .alu_out_Q103H(alu_out_Q103H),
    .dmem_wr_data_Q103H(dmem_wr_data_Q103H),
    .dmem_wr_en_Q103H(dmem_wr_en_Q103H),
    .dmem_byte_en_Q103H(dmem_byte_en_Q103H),
    .dmem_is_signed_Q103H(dmem_is_signed_Q103H),
    .dmem_rd_data_Q104H(dmem_rd_data_Q104H)
  );

  // ============================
  // Instruction memory image
  // ============================
  logic [31:0] IMem [0:IMEM_SIZE_WORDS-1];

  initial begin
    clk = 0;
    rst = 1;
    ready_Q101H = 0;

    pc_Q100H = 0;
    alu_out_Q103H = 0;
    dmem_wr_data_Q103H = 0;
    dmem_wr_en_Q103H = 0;
    dmem_byte_en_Q103H = 4'b1111;
    dmem_is_signed_Q103H = 0;

    // ==========================================================
    // FIXED: Load instruction memory directly via hierarchy
    // No 'force' statement needed.
    // Assuming the array inside d_mem is named 'mem'.
    // ==========================================================
    $display("TB: Loading instruction memory directly into DUT");
    $readmemh("verif/memory/inst_mem.hex", dut.i_mem.mem);


    // ============================
    // Load instruction memory
    // ============================
    //$display("TB: Loading instruction memory using readmemh");
    //$readmemh("inst_mem.hex", IMem);

    // ============================
    // Backdoor force into I_MEM
    // ============================
    //$display("TB: Forcing IMem into DUT instruction memory");
    //force dut.i_mem.mem = IMem;

    #20;
    rst = 0;
    ready_Q101H = 1;

    // ============================
    // Fetch few instructions
    // ============================
    repeat (5) begin
      @(posedge clk);
      $display("PC=0x%08h -> INSTR=0x%08h",
               pc_Q100H, instruction_Q101H);
      pc_Q100H += 4;
    end

    // ============================
    // Data memory write
    // ============================
    $display("TB: Writing to D_MEM");
    @(posedge clk);
    alu_out_Q103H = 32'h00000010;
    dmem_wr_data_Q103H = 32'hDEADBEEF;
    dmem_wr_en_Q103H = 1;

    @(posedge clk);
    dmem_wr_en_Q103H = 0;

    // ============================
    // Data memory read
    // ============================
    @(posedge clk);
    alu_out_Q103H = 32'h00000010;

    @(posedge clk);
    $display("D_MEM READ DATA = 0x%08h", dmem_rd_data_Q104H);

    // ============================
    // Finish
    // ============================
    $display("TB: Finished successfully");
    #20;
    $finish;
  end

endmodule
